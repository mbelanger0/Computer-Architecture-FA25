`include "memory.sv"
`include "ws2812b.sv"
`include "controller.sv"

// led_matrix top level module

module top(
    input logic     clk, 
    input logic     SW, 
    input logic     BOOT, 
    output logic    _48b, 
    output logic    _45a
);

    logic [7:0] red_data;
    logic [7:0] green_data;
    logic [7:0] blue_data;

    logic [5:0] pixel;
    logic [4:0] frame;
    logic [10:0] address;

    logic [23:0] shift_reg = 24'd0;
    logic load_sreg;
    logic transmit_pixel;
    logic shift;
    logic ws2812b_out;

    assign address = { frame, pixel };

    // Instance sample memory for red channel
    memory #(
        .INIT_FILE      ("spiral/red.txt")
    ) u1 (
        .clk            (clk), 
        .read_address   (address), 
        .read_data      (red_data)
    );

    // Instance sample memory for green channel
    memory #(
        .INIT_FILE      ("spiral/green.txt")
    ) u2 (
        .clk            (clk), 
        .read_address   (address), 
        .read_data      (green_data)
    );

    // Instance sample memory for blue channel
    memory #(
        .INIT_FILE      ("spiral/blue.txt")
    ) u3 (
        .clk            (clk), 
        .read_address   (address), 
        .read_data      (blue_data)
    );

    // Instance the WS2812B output driver
    ws2812b u4 (
        .clk            (clk), 
        .serial_in      (shift_reg[23]), 
        .transmit       (transmit_pixel), 
        .ws2812b_out    (ws2812b_out), 
        .shift          (shift)
    );

    // Instance the controller
    controller u5 (
        .clk            (clk), 
        .load_sreg      (load_sreg), 
        .transmit_pixel (transmit_pixel), 
        .pixel          (pixel), 
        .frame          (frame)
    );

    // // ***LEDs flashing for testing and debugging***
    
    // parameter FLASH_INTERVAL = 6000000;
    // logic [$clog2(FLASH_INTERVAL) - 1:0] count = 0;
    // logic flash_on = 1'b0;

    // always_ff @(posedge clk) begin
    //     if (count == FLASH_INTERVAL - 1) begin
    //         count <= 0;
    //         flash_on <= ~flash_on;
    //     end else begin
    //         count <= count + 1;
    //     end

    //     if (load_sreg) begin
    //         shift_reg <= flash_on ? 24'h080808 : 24'h000000;
    //     end else if (shift) begin
    //         shift_reg <= { shift_reg[22:0], 1'b0 };
    //     end
    // end
            
    

    always_ff @(posedge clk) begin
        if (load_sreg) begin
            unique case ({ SW, BOOT })
                2'b00:
                    shift_reg <= { green_data, 16'd0 };
                2'b01:
                    shift_reg <= { 8'd0, red_data, 8'd0 };
                2'b10:
                    shift_reg <= { 16'd0, blue_data };
                2'b11:
                    shift_reg <= { green_data, red_data, blue_data };
            endcase
        end
        else if (shift) begin
            shift_reg <= { shift_reg[22:0], 1'b0 };
        end
    end

    assign _48b = ws2812b_out;
    assign _45a = ~ws2812b_out;

endmodule
